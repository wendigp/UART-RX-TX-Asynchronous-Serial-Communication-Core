
module baud_rate_gen_rx #(
			parameter CLK_FREQ = 50_000_000,
			parameter BAUD_RATE = 9600)(
			input wire clk,
			input wire rst_n,
			output reg sample_tick);		//16x baud tick

localparam integer SAMPLE_MAX_CNT = CLK_FREQ / (BAUD_RATE * 16);
reg [$clog2(SAMPLE_MAX_CNT)-1 : 0] sample_cnt;

always @(posedge clk, negedge rst_n)
begin
	if(!rst_n)
		begin
		sample_tick <= 1'b0;
		sample_cnt  <= 0;
		end
	else
		begin
			if(sample_cnt == SAMPLE_MAX_CNT)
				begin
				sample_tick <= 1'b1;
				sample_cnt <= 0;
				end
			else
				begin
				sample_tick <= 1'b0;
				sample_cnt <= sample_cnt + 1;
				end
		end
end
endmodule
