//TB

module uart_tb;
	
//CLOCK & RESET
	reg clk;
	reg rst_n;
	
//TX INTERFACE
	reg [7:0]tx_data;
	reg tx_start;
	wire tx_busy;
	wire tx_serial;

//RX INTERFACE
	wire [7:0]rx_data;
	wire data_ready;

//DUT 
uart_top DUT(
		.clk(clk),
		.reset_n(rst_n),
		.tx_start(tx_start),
		.tx_data(tx_data),
		.tx_busy(tx_busy),
		.tx_serial(tx_serial),

		.rx_serial(tx_serial),
		.rx_data(rx_data),
		.data_ready(data_ready)
		);

//===============CLOCK GEN - 50MHz===============//
initial
clk = 0;
always #10 clk = ~clk;

//=================RESET========================//
initial
	begin
	rst_n = 0;
	tx_start = 0;
	tx_data = 8'd0;
	#200;
	rst_n = 1;
	end

task send_byte (input [7:0]data);
	begin
	while(tx_busy)
		@(posedge clk)

	@(posedge clk)
	tx_data <= data;
	tx_start <= 1'b1;

	@(posedge clk)
	tx_start <= 1'b0;
	end
endtask

//TEST SEQUENCE
  initial begin
    @(posedge rst_n);

 // Test 1
    send_byte(8'h55);
    wait(data_ready);
    if (rx_data !== 8'h55)
      $display("? ERROR: Expected 55, got %h", rx_data);
    else
      $display("? PASS: 55");

    // Test 2
    send_byte(8'hA3);
    wait(data_ready)
    if (rx_data !== 8'hA3)
      $display("? ERROR: Expected A3, got %h", rx_data);
    else
      $display("? PASS: A3");

 // Test 3
    send_byte(8'hFF);
    wait(data_ready)
    if (rx_data !== 8'hFF)
      $display("? ERROR: Expected FF, got %h", rx_data);
    else
      $display("? PASS: FF");

    $display("?? UART LOOPBACK TEST COMPLETED SUCCESSFULLY");
    #1000;
    $stop;
  end

endmodule
		
